`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2021/04/04 17:00:56
// Design Name:
// Module Name: FA
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module FA(a, b, c_in, s, c_out);
  input a,b,c_in;
  output s,c_out;
  
  assign s = a^b^c_in;
  assign c_out=(a&b)|(b&c_in)|(c_in&a);
  
endmodule
